library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mouse_hunt is
    port (
        
    );
end entity mouse_hunt;

architecture rtl of mouse_hunt is
    
    component mouse_hunt_fd is
        port (
            
        );
    end component;

    component mouse_hunt_uc is
        port (
            
        );
    end component;

begin
    
    
    
end architecture rtl;