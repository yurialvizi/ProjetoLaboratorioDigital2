library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mouse_hunt_uc is
    port (
        
    );
end entity mouse_hunt_uc;

architecture rtl of mouse_hunt_uc is
    
begin
    
    
    
end architecture rtl;